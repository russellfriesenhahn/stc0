`define CMDADDRH                            31
`define CMDADDRL                            8
`define CMDH                                7
`define CMDL                                0
`define CTRLWRD_SZ                          10
`define CTRL_BF0                            0
`define CTRL_ES                             13
`define LASTWORD                            16'habcd
`define RAH                                 5
`define RAL                                 2
`define RA_BFP_CTRL0                        8'h00
`define RA_BFP_STAT0                        8'h04
`define RA_CTRL_BFP                         4'ha
`define RA_CTRL_CTRL0                       4'h0
`define RA_CTRL_CTRL1                       4'h1
`define RA_CTRL_CTRLWORD                    7
`define RA_CTRL_LFSRS_CTRL                  2
`define RA_CTRL_LFSRS_ITERATIONS            4
`define RA_CTRL_LFSRS_STRIDE                3
`define RA_CTRL_LFSRX_SEED                  5
`define RA_CTRL_LFSRY_SEED                  6
`define RA_CTRL_MUXCTRL                     8'h01
`define RA_CTRL_STAT0                       4'h2
`define RA_CTRL_STAT1                       4'h3
`define RA_CTRL_XINGRESS                    4'h8
`define RA_CTRL_YINGRESS                    4'h9
`define RB_BFCTRL_BFBYPASS                  4
`define RB_BFCTRL_BFBYPASSX                 5
`define RB_BFCTRL_SS                        0
`define RB_BFCTRL_TWRD                      6
`define RB_BFCTRL_TWWR                      7
`define RB_CTRL_ADDR                        28
`define RB_EGRESSCTRL_CRCBYPASS             3
`define RB_EGRESSCTRL_OUTPUTEN              2
`define RB_EGRESSCTRL_OUTPUTMUX             0
`define RB_LFSRCTRL_ENABLE                  0
`define RB_LFSRCTRL_ITERS                   65536
`define RB_LFSRCTRL_ITERSRC                 1
`define RB_LFSRCTRL_STRIDE                  256
`define RMH                                 21
`define RML                                 14
`define RM_CTRL                             8'h01
`define RM_XYINGRESS                        8'h03
`define WRITE                               8'h01
